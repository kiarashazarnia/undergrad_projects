module Adder12(
    input [11:0]a,b,
    output [11:0] w);
    assign w = a + b;
endmodule