module InsMemory (
	input[11:0]  address,
	output[18:0]  ins_out
);
	logic[18:0] ins [4095:0];
    initial begin
		/*case 1*/
        // 	 ins[0] = 19'b1000000100001100100;
		//  ins[1] = 19'b1000001000001100110;
		//  ins[2] = 19'b0000001100101000000;
		//  ins[3] = 19'b1000101100001101000;
		//  ins[4] = 19'b1000000100001100101;
		//  ins[5] = 19'b1000001000001100111;
		//  ins[6] = 19'b0000101100101000000;
		//  ins[7] = 19'b1000101100001101001;
		/*case 2*/
		ins[0] = 19'b0000011100000000000;
		ins[1] = 19'b0000000100000000000;
		ins[2] = 19'b0101001100100010100;
		ins[3] = 19'b1010000000000001010;//4+?6DISP + PC+1
		ins[4] = 19'b1000001000101100100;
		ins[5] = 19'b0001001111101000000;
		ins[6] = 19'b1011100000000000001;
		ins[7] = 19'b0000011101000000000;
		ins[8] = 19'b0100000100100000001;
		ins[9] = 19'b1110000000000000010;
    end
	assign ins_out = ins[address];
endmodule
