module PCAdd1(
	input[11:0]  pcIn,
	output[11:0] pcOut
);
	assign pcOut = pcIn + 1;
endmodule


